`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name: lab1
//////////////////////////////////////////////////////////////////////////////////


module counter(clk, out);
input clk;                    // ����ʱ��
output [2:0] out;             // ����ֵ

always @(posedge clk)  begin  // ��ʱ�������ؼ�������1
    out <= out + 1;                        // ����ʵ��
end                           
endmodule



