`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name: lab1
//////////////////////////////////////////////////////////////////////////////////


module dynamic _scan(clk,  SEG, AN);
input clk;              // ϵͳʱ��
output [7:0] SEG;  		// �ֱ��ӦCA��CB��CC��CD��CE��CF��CG��DP
output [7:0] AN;        // 8λ�����Ƭѡ�ź�
assign AN[7:0] = 
                      // ����ʵ��
endmodule



